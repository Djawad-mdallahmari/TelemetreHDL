module Compteur(clk,signalCapteur,cnt);

input clk,signalCapteur;
output reg[15:0] cnt;

always@(negedge(clk))
begin
	if(signalCapteur)
	begin
		cnt <= cnt + 1;
	end
	else
	begin
		cnt <= 0;
	end
end

endmodule
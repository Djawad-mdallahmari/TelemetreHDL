module Telemetre(CLOCK_50,SMA_CLKIN,HEX0,HEX1,HEX2,LEDR6);

input CLOCK_50,SMA_CLKIN;
output reg[7:0] HEX0,HEX1,HEX2;
output LEDR6;


endmodule